library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity testALU is
end entity;

architecture test of testALU is
  component ArithmeticUnit is
    port (
    A : in std_logic_vector(15 downto 0);
    B : in std_logic_vector(15 downto 0);
    --  B -> Rs   and A -> RD
    funcSelect : in std_logic_vector(3 downto 0);
    -- funcSelect is considered with optional parts  TODO : handle optionals later
    Cin  : in std_logic;
    Zin  : in std_logic;
    Cout  : out std_logic;
    Zout  : out std_logic;
    --  z  is Zeroflag
    AluOut_on_Databus : out std_logic_vector(15 downto 0) 
    );
end component;

  signal A : std_logic_vector (15 downto 0);
  signal B : std_logic_vector (15 downto 0);
  signal funcSelect : std_logic_vector(3 downto 0);
  signal Cin : std_logic;
  signal Zin : std_logic;
  signal Cout : std_logic;
  signal Zout : std_logic;
  signal AluOut_on_Databus : std_logic_vector(15 downto 0);

  begin
    an : ArithmeticUnit port map (A => A , B => B , funcSelect => funcSelect , Cin => Cin , Zin => Zin , Cout => Cout, Zout => Zout ,AluOut_on_Databus => AluOut_on_Databus);
    A <= "1101101001011100";
    B <= "0010111000101101";
    funcSelect <= "1001";--,"0001" after 100 ns , "0010" after 200 ns , "0011" after 300 ns , "0100" after 400 ns , "0101" after 510 ns , "0110" after 600 ns , "0111" after 700 ns , "1000" after 800 ns;
    Cin <= '0';
    Zin <= '0';
end test;